library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ALUControl is
	port(ALUOp : in std_logic_vector(1 downto 0);
			functCode : in std_logic_vector(5 downto 0);
			ALUCont : out std_logic_vector(3 downto 0));
end ALUControl;

architecture control of ALUControl is
begin
process(ALUOp,functCode)
begin
	case ALUOp is
		when "00" => ALUCont <= "0010";
		when "01" => ALUCont <= "0110";
		when "10" =>
			case functCode is
				when "100000" => ALUCont <= "0010";
				when "100010" => ALUCont <= "0110";
				when "100100" => ALUCont <= "0000";
				when "100101" => ALUCont <= "0001";
				when "101010" => ALUCont <= "0111";
				when "100111" => ALUCont <= "1100";
				when others => ALUCont <= "0000";
			end case;
		when others => ALUCont <= "0000";
	end case;
end process;
end control;