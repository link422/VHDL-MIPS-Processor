library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity decoder is
port( x : in std_logic_vector (4 downto 0);
		regNum : out std_logic_vector (31 downto 0));
end decoder;

architecture decode of decoder is
begin
process(x)
begin
	case x is 
		when "00000" => regNum <= "00000000000000000000000000000001";
		when "00001" => regNum <= "00000000000000000000000000000010";
		when "00010" => regNum <= "00000000000000000000000000000100";
		when "00011" => regNum <= "00000000000000000000000000001000";
		when "00100" => regNum <= "00000000000000000000000000010000";
		when "00101" => regNum <= "00000000000000000000000000100000";
		when "00110" => regNum <= "00000000000000000000000001000000";
		when "00111" => regNum <= "00000000000000000000000010000000";
		when "01000" => regNum <= "00000000000000000000000100000000";
		when "01001" => regNum <= "00000000000000000000001000000000";
		when "01010" => regNum <= "00000000000000000000010000000000";
		when "01011" => regNum <= "00000000000000000000100000000000";
		when "01100" => regNum <= "00000000000000000001000000000000";
		when "01101" => regNum <= "00000000000000000010000000000000";
		when "01110" => regNum <= "00000000000000000100000000000000";
		when "01111" => regNum <= "00000000000000001000000000000000";
		when "10000" => regNum <= "00000000000000010000000000000000";
		when "10001" => regNum <= "00000000000000100000000000000000";
		when "10010" => regNum <= "00000000000001000000000000000000";
		when "10011" => regNum <= "00000000000010000000000000000000";
		when "10100" => regNum <= "00000000000100000000000000000000";
		when "10101" => regNum <= "00000000001000000000000000000000";
		when "10110" => regNum <= "00000000010000000000000000000000";
		when "10111" => regNum <= "00000000100000000000000000000000";
		when "11000" => regNum <= "00000001000000000000000000000000";
		when "11001" => regNum <= "00000010000000000000000000000000";
		when "11010" => regNum <= "00000100000000000000000000000000";
		when "11011" => regNum <= "00001000000000000000000000000000";
		when "11100" => regNum <= "00010000000000000000000000000000";
		when "11101" => regNum <= "00100000000000000000000000000000";
		when "11110" => regNum <= "01000000000000000000000000000000";
		when "11111" => regNum <= "10000000000000000000000000000000";
		when others  => regNum <= "00000000000000000000000000000000";
	end case;
end process;
end decode;
		
