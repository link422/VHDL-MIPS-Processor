library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity signExtend is
port (in1 : in std_logic_vector (15 downto 0);
		out1 : out std_logic_vector (31 downto 0));
end signExtend;

architecture arch of signExtend is
signal temp : std_logic_vector (31 downto 0);
begin
process(in1)
begin
	IF in1(15) = '1' THEN
		temp(31 downto 16) <= "1111111111111111";
	ELSE
		temp(31 downto 16) <= "0000000000000000";
	END IF;
	temp(15 downto 0) <= in1;
		
end process;
out1 <= temp;
end arch;