library ieee;
use ieee.std_logic_1164.all;

package multiplex_pack is
        type regArray is array(31 downto 0) of std_logic_vector (31 downto 0);
end package;