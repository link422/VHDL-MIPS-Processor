library ieee;
use ieee.std_logic_1164.all;

entity sevSeg is
	port(x : in std_logic_vector(7 downto 0);
			o1,o2 : out std_logic_vector(7 downto 0));
end sevSeg;

architecture sev of sevSeg is
begin
process(x)
begin
	case x is
		when "00000000" =>   --00
			o1 <= "11000000";
			o2 <= "11000000";
		when "00000001" =>	--01
			o1 <= "11111001";
			o2 <= "11000000";
		when "00000010" =>	--02
			o1 <= "10100100";
			o2 <= "11000000";
		when "00000011" =>	--03
			o1 <= "10110000";
			o2 <= "11000000";
		when "00000100" =>	--04
			o1 <= "10011001";
			o2 <= "11000000";
		when "00000101" =>	--05
			o1 <= "10010010";
			o2 <= "11000000";
		when "00000110" =>	--06
			o1 <= "10000010";
			o2 <= "11000000";
		when "00000111" =>	--07
			o1 <= "11111000";
			o2 <= "11000000";
		when "00001000" =>	--08
			o1 <= "10000000";
			o2 <= "11000000";
		when "00001001" =>	--09
			o1 <= "10010000";
			o2 <= "11000000";
		when "00001010" =>	--0a
			o1 <= "10100000";
			o2 <= "11000000";
		when "00001011" =>	--0b
			o1 <= "10000011";
			o2 <= "11000000";
		when "00001100" =>	--0c
			o1 <= "10100111";
			o2 <= "11000000";
		when "00001101" =>	--0d
			o1 <= "10100001";
			o2 <= "11000000";
		when "00001110" =>	--0e
			o1 <= "10000110";
			o2 <= "11000000";
		when "00001111" =>	--0f
			o1 <= "10001110";
			o2 <= "11000000";
		when "00010000" =>   --10
			o1 <= "11000000";
			o2 <= "11111001";
		when "00010001" =>	--11
			o1 <= "11111001";
			o2 <= "11111001";
		when "00010010" =>	--12
			o1 <= "10100100";
			o2 <= "11111001";
		when "00010011" =>	--13
			o1 <= "10110000";
			o2 <= "11111001";
		when "00010100" =>	--14
			o1 <= "10011001";
			o2 <= "11111001";
		when "00010101" =>	--15
			o1 <= "10010010";
			o2 <= "11111001";
		when "00010110" =>	--16
			o1 <= "10000010";
			o2 <= "11111001";
		when "00010111" =>	--17
			o1 <= "11111000";
			o2 <= "11111001";
		when "00011000" =>	--18
			o1 <= "10000000";
			o2 <= "11111001";
		when "00011001" =>	--19
			o1 <= "10010000";
			o2 <= "11111001";
		when "00011010" =>	--1a
			o1 <= "10100000";
			o2 <= "11111001";
		when "00011011" =>	--1b
			o1 <= "10000011";
			o2 <= "11000000";
		when "00011100" =>	--1c
			o1 <= "10100111";
			o2 <= "11111001";
		when "00011101" =>	--1d
			o1 <= "10100001";
			o2 <= "11111001";
		when "00011110" =>	--1e
			o1 <= "10000110";
			o2 <= "11111001";
		when "00011111" =>	--1f
			o1 <= "10001110";
			o2 <= "11111001";
		when "00101111" =>	--2f
			o1 <= "10001110";
			o2 <= "10100100";
		when "00111111" =>	--3f
			o1 <= "10001110";
			o2 <= "10110000";
		when "01001111" =>	--4f
			o1 <= "10001110";
			o2 <= "10011001";
		when "01011111" =>	--5f
			o1 <= "10001110";
			o2 <= "10010010";
		when "01101111" =>	--6f
			o1 <= "10001110";
			o2 <= "10000010";
		when "01111111" =>	--7f
			o1 <= "10001110";
			o2 <= "11111000";
		when "10001111" =>	--8f
			o1 <= "10001110";
			o2 <= "10000000";
		when "10011111" =>	--9f
			o1 <= "10001110";
			o2 <= "10010000";
		when "10101111" =>	--af
			o1 <= "10001110";
			o2 <= "10100000";
		when "10111111" =>	--bf
			o1 <= "10001110";
			o2 <= "10000011";
		when "11001111" =>	--cf
			o1 <= "10001110";
			o2 <= "10100111";
		when "11011111" =>	--df
			o1 <= "10001110";
			o2 <= "10100001";
		when "11101111" =>	--ef
			o1 <= "10001110";
			o2 <= "10000110";
		when "11111111" =>	--ff
			o1 <= "10001110";
			o2 <= "10001110";
		when others =>
			o1 <= "--------";
			o2 <= "--------";
	end case;
end process;
end sev;