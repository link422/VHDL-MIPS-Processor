library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity add_block is
port (in1 : in std_logic_vector (31 downto 0);
		in2 : in std_logic_vector (31 downto 0);
		out1 : out std_logic_vector (31 downto 0));
end add_block;

architecture add of add_block is
signal temp : std_logic_vector (31 downto 0);
begin
process(in1)
begin
	temp <= in1 + in2;
end process;
out1 <= temp;
end add;